// outline for the module:
// use cordic to calculate the I and the Q values of the input with just
// a zero value at the input y of the incoming cordic module
// 
